VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_power_routing
  CLASS BLOCK ;
  FOREIGN caravel_power_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
END caravel_power_routing



END LIBRARY

