VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_signal_routing
  CLASS BLOCK ;
  FOREIGN caravan_signal_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;


END caravan_signal_routing
END LIBRARY

